entity E1 is
port(A: in natural:=1;
B:inout natural:=1);
end ent